// Implements Nios II system for the DE1-SoC Board
// Inputs:  SW7-0 are parallel port inputs to the Nios II system
//          CLOCK_50 is the system clock (50MHz)
//          KEY0 is the active-low system reset
// Outputs: LEDR7-0 are parallel port outputs from the Nios II system

module task4(CLOCK_50, SW, KEY, LEDR,
             VGA_R, VGA_G, VGA_B,
             VGA_HS, VGA_VS, VGA_CLK);

  input CLOCK_50;
  input [7:0] SW;
  input [3:0] KEY;
  output [7:0] LEDR;

  output [7:0] VGA_R, VGA_G, VGA_B;
  output VGA_HS, VGA_VS, VGA_CLK;

  // Instantiate NiosII system module generated by the Qsys Tool
  pixel_xform_system u0 (
      .clk_clk         (CLOCK_50),    // clk.clk
      .leds_export     (LEDR),        // leds.export
      .reset_reset_n   (KEY[0]),      // reset.reset_n
      .switches_export (SW),          // switches.export
      .vga_b_readdata               (VGA_B),
      .vga_clk_writeresponsevalid_n (VGA_CLK),
      .vga_g_readdata               (VGA_G),
      .vga_hs_writeresponsevalid_n  (VGA_HS),
      .vga_r_readdata               (VGA_R),
      .vga_vs_writeresponsevalid_n  (VGA_VS)
  );

endmodule
