// Implements Nios II system for the DE1-SoC Board
// Inputs:  SW7-0 are parallel port inputs to the Nios II system
//          CLOCK_50 is the system clock (50MHz)
//          KEY0 is the active-low system reset
// Outputs: LEDR7-0 are parallel port outputs from the Nios II system

module task2(CLOCK_50, SW, KEY, LEDR);

  input CLOCK_50;
  input [7:0] SW;
  input [3:0] KEY;
  output [7:0] LEDR;

  // Instantiate NiosII system module generated by the Qsys Tool
  pixel_xform_system u0 (
      .clk_clk         (CLOCK_50),    // clk.clk
      .leds_export     (LEDR),        // leds.export
      .reset_reset_n   (KEY[0]),      // reset.reset_n
      .switches_export (SW)           // switches.export
  );

endmodule
